module moore_model
