module MEMORY_CELL(
  input select,
  input read_write,
  input in,
  output reg out
);
endmodule
