module NOT_GATE (input a, output y);
  assign y = ~a;
endmodule
