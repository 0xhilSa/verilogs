module WAVE (
  input wire wave
);
endmodule
